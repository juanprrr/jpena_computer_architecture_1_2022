/* 
	Instruction Memory.
	Set Default ARM Instructions
*/

module instructionMemory(input logic[7:0] address, //Memory Address in range [0-255] -> 2^8
								 output logic[16:0] data	  //Read data value -> read value port 
								 );
	always @*
		case(address)
				17b'00000000000000000: data = 17b'00001111011111111;
				17b'00000000000000100: data = 17b'00100111000100010;
				17b'00000000000001000: data = 17b'00100111000010111;
				17b'00000000000001100: data = 17b'01000001000010000;
				17b'00000000000010000: data = 17b'01001010000010000;
				17b'00000000000010100: data = 17b'00000010101000010;
				17b'00000000000011000: data = 17b'10000000000000001;
				17b'00000000000011100: data = 17b'00010001011110100;
				17b'00000000000100000: data = 17b'10000011111111111;
				17b'00000000000100100: data = 17b'00000111010000010;
				17b'00000000000101000: data = 17b'00000111010000010;
				17b'00000000000101100: data = 17b'00000000000000000;
				17b'00000000000110000: data = 17b'00000000000000000:
			
			default: data = 17'b0;
			
			
		endcase 

endmodule